magic
tech scmos
timestamp 1731099534
<< nwell >>
rect -33 -13 38 70
<< polysilicon >>
rect -20 46 -19 50
rect 20 47 21 51
rect -20 43 -18 46
rect 20 43 22 47
rect -20 -7 -18 -1
rect 20 -6 22 -1
rect -20 -28 -18 -23
rect 20 -28 22 -23
rect -20 -35 -18 -33
rect 20 -35 22 -33
rect -20 -39 -19 -35
rect 20 -39 21 -35
<< ndiffusion >>
rect -25 -29 -20 -28
rect -22 -33 -20 -29
rect -18 -32 -17 -28
rect -18 -33 -13 -32
rect 19 -32 20 -28
rect 15 -33 20 -32
rect 22 -32 23 -28
rect 22 -33 27 -32
<< pdiffusion >>
rect -21 39 -20 43
rect -25 31 -20 39
rect -21 27 -20 31
rect -25 17 -20 27
rect -21 13 -20 17
rect -25 3 -20 13
rect -21 -1 -20 3
rect -18 39 -17 43
rect -18 31 -13 39
rect -18 27 -17 31
rect -18 17 -13 27
rect -18 13 -17 17
rect -18 3 -13 13
rect -18 -1 -17 3
rect 19 39 20 43
rect 15 31 20 39
rect 19 27 20 31
rect 15 17 20 27
rect 19 13 20 17
rect 15 3 20 13
rect 19 -1 20 3
rect 22 39 23 43
rect 22 31 27 39
rect 22 27 23 31
rect 22 17 27 27
rect 22 13 23 17
rect 22 3 27 13
rect 22 -1 23 3
<< metal1 >>
rect -32 67 34 68
rect -32 63 -26 67
rect -22 63 -11 67
rect -7 63 7 67
rect 11 63 24 67
rect 28 63 34 67
rect -32 62 34 63
rect -25 43 -22 62
rect -15 46 -11 50
rect 25 47 29 51
rect -13 39 15 43
rect 23 -28 27 -1
rect -13 -32 15 -28
rect -26 -47 -22 -33
rect -15 -39 -11 -35
rect 25 -39 29 -35
rect -34 -48 38 -47
rect -34 -52 -26 -48
rect -22 -52 -8 -48
rect -4 -52 8 -48
rect 12 -52 24 -48
rect 28 -52 38 -48
rect -34 -53 38 -52
<< ntransistor >>
rect -20 -33 -18 -28
rect 20 -33 22 -28
<< ptransistor >>
rect -20 -1 -18 43
rect 20 -1 22 43
<< polycontact >>
rect -19 46 -15 50
rect 21 47 25 51
rect -19 -39 -15 -35
rect 21 -39 25 -35
<< ndcontact >>
rect -26 -33 -22 -29
rect -17 -32 -13 -28
rect 15 -32 19 -28
rect 23 -32 27 -28
<< pdcontact >>
rect -25 39 -21 43
rect -25 27 -21 31
rect -25 13 -21 17
rect -25 -1 -21 3
rect -17 39 -13 43
rect -17 27 -13 31
rect -17 13 -13 17
rect -17 -1 -13 3
rect 15 39 19 43
rect 15 27 19 31
rect 15 13 19 17
rect 15 -1 19 3
rect 23 39 27 43
rect 23 27 27 31
rect 23 13 27 17
rect 23 -1 27 3
<< psubstratepcontact >>
rect -26 -52 -22 -48
rect -8 -52 -4 -48
rect 8 -52 12 -48
rect 24 -52 28 -48
<< nsubstratencontact >>
rect -26 63 -22 67
rect -11 63 -7 67
rect 7 63 11 67
rect 24 63 28 67
<< labels >>
rlabel metal1 -13 48 -13 48 1 Vbias1
rlabel metal1 -1 65 -1 65 5 Vdd
rlabel metal1 27 49 27 49 1 Vbias2
rlabel metal1 -13 -37 -13 -37 1 Vin
rlabel metal1 27 -37 27 -37 1 Vbias3
rlabel metal1 1 -50 1 -50 1 GND
rlabel metal1 27 -19 27 -17 1 Vout
<< end >>
