magic
tech scmos
timestamp 1699311399
<< nwell >>
rect -46 283 88 336
rect 66 282 78 283
<< ntransistor >>
rect -29 248 -27 253
rect -7 243 -5 253
rect 15 243 17 253
rect 37 243 39 253
rect -7 201 -5 211
rect 15 201 17 211
rect 37 201 39 211
<< ptransistor >>
rect -29 294 -27 318
rect -7 294 -5 318
rect 15 310 17 318
rect 37 294 39 318
rect 59 294 61 318
<< ndiffusion >>
rect -34 252 -29 253
rect -31 248 -29 252
rect -27 252 -26 253
rect -27 249 -22 252
rect -27 248 -26 249
rect -12 247 -7 253
rect -8 243 -7 247
rect -5 249 -4 253
rect -5 243 0 249
rect 10 250 15 253
rect 14 246 15 250
rect 10 243 15 246
rect 17 249 20 253
rect 32 250 37 253
rect 17 243 22 249
rect 36 246 37 250
rect 32 243 37 246
rect 39 249 40 253
rect 39 243 44 249
rect -14 208 -7 211
rect -10 204 -7 208
rect -14 201 -7 204
rect -5 209 0 211
rect -5 205 -4 209
rect -5 201 0 205
rect 10 208 15 211
rect 14 204 15 208
rect 10 201 15 204
rect 17 209 22 211
rect 17 205 18 209
rect 17 201 22 205
rect 32 208 37 211
rect 36 204 37 208
rect 32 201 37 204
rect 39 209 44 211
rect 39 205 40 209
rect 39 201 44 205
<< pdiffusion >>
rect -30 314 -29 318
rect -34 294 -29 314
rect -27 303 -22 318
rect -27 299 -26 303
rect -27 294 -22 299
rect -8 314 -7 318
rect -12 294 -7 314
rect -5 314 -1 318
rect 14 314 15 318
rect -5 303 0 314
rect 10 310 15 314
rect 17 314 24 318
rect 17 310 20 314
rect 36 314 37 318
rect -5 299 -4 303
rect -5 294 0 299
rect 32 294 37 314
rect 39 303 44 318
rect 39 299 40 303
rect 39 294 44 299
rect 58 314 59 318
rect 54 294 59 314
rect 61 302 66 318
rect 61 298 62 302
rect 61 294 66 298
<< ndcontact >>
rect -35 248 -31 252
rect -26 252 -22 256
rect -26 245 -22 249
rect -12 243 -8 247
rect -4 249 0 253
rect 10 246 14 250
rect 20 249 24 253
rect 32 246 36 250
rect 40 249 44 253
rect -14 204 -10 208
rect -4 205 0 209
rect 10 204 14 208
rect 18 205 22 209
rect 32 204 36 208
rect 40 205 44 209
<< pdcontact >>
rect -34 314 -30 318
rect -26 299 -22 303
rect -12 314 -8 318
rect -1 314 3 318
rect 10 314 14 318
rect 20 310 24 314
rect 32 314 36 318
rect -4 299 0 303
rect 40 299 44 303
rect 54 314 58 318
rect 62 298 66 302
<< nsubstratencontact >>
rect -34 327 -30 331
rect -12 327 -8 331
rect 10 327 14 331
rect 32 327 36 331
rect 50 327 54 331
<< polysilicon >>
rect -29 318 -27 324
rect -7 318 -5 324
rect 15 318 17 324
rect 59 321 60 325
rect 37 318 39 321
rect 59 318 61 321
rect 15 307 17 310
rect 15 300 17 303
rect -29 292 -27 294
rect -7 292 -5 294
rect 37 292 39 294
rect 59 292 61 294
rect -29 288 -28 292
rect -6 288 -5 292
rect 38 288 39 292
rect 60 288 61 292
rect -29 284 -27 288
rect -28 280 -27 284
rect -29 253 -27 260
rect -7 253 -5 260
rect 15 253 17 260
rect 37 253 39 260
rect -29 241 -27 248
rect -29 237 -28 241
rect -7 233 -5 243
rect 15 239 17 243
rect 15 237 16 239
rect 37 237 39 243
rect -7 217 -5 220
rect 16 217 17 221
rect -6 213 -5 217
rect -7 211 -5 213
rect 15 211 17 217
rect 37 211 39 217
rect -7 195 -5 201
rect 15 195 17 201
rect 37 195 39 201
rect -7 191 -6 195
rect 15 191 16 195
rect 37 191 38 195
<< polycontact >>
rect 60 321 64 325
rect 13 303 17 307
rect 15 296 19 300
rect -28 288 -24 292
rect -10 288 -6 292
rect 34 288 38 292
rect 56 288 60 292
rect -32 280 -28 284
rect -31 260 -27 264
rect -8 260 -4 264
rect 14 260 18 264
rect 35 260 39 264
rect -28 237 -24 241
rect 16 235 20 239
rect 12 217 16 221
rect -10 213 -6 217
rect -6 191 -2 195
rect 16 191 20 195
rect 38 191 42 195
<< metal1 >>
rect -37 331 66 333
rect -37 327 -34 331
rect -30 327 -12 331
rect -8 327 10 331
rect 14 327 32 331
rect 36 327 50 331
rect 54 328 66 331
rect -34 318 -30 327
rect -12 318 -8 327
rect 10 318 14 327
rect 54 318 57 328
rect 44 299 45 302
rect 15 292 19 296
rect -24 288 -10 292
rect 15 288 34 292
rect -37 280 -32 284
rect 28 279 32 288
rect 41 271 45 299
rect 60 288 62 291
rect 58 271 62 288
rect 41 268 62 271
rect -27 260 -8 264
rect -4 260 14 264
rect 18 260 35 264
rect 58 253 62 268
rect -26 241 -22 245
rect -24 237 -22 241
rect -15 243 -12 247
rect 44 249 62 253
rect -15 229 -11 243
rect 10 229 13 246
rect 32 229 36 246
rect -15 225 0 229
rect 10 225 22 229
rect 32 225 44 229
rect -3 209 0 225
rect 19 209 22 225
rect 40 209 44 225
rect -2 191 16 195
rect 20 191 38 195
rect -39 186 64 187
rect -39 185 10 186
rect -39 180 -34 185
rect -29 180 -14 185
rect -9 181 10 185
rect 15 181 32 186
rect 37 181 64 186
rect -9 180 64 181
rect -39 178 64 180
<< m2contact >>
rect -34 180 -29 185
rect -14 180 -9 185
rect 10 181 15 186
rect 32 181 37 186
<< metal2 >>
rect 32 322 51 326
rect -4 314 7 318
rect 32 314 36 322
rect -26 252 -22 303
rect -34 185 -30 251
rect -4 249 0 303
rect 4 217 7 314
rect 20 307 24 314
rect 13 303 24 307
rect 20 249 24 303
rect 47 286 51 322
rect 60 321 69 325
rect 62 286 66 302
rect 47 282 66 286
rect 16 235 23 239
rect 13 217 25 221
rect -9 213 7 217
rect -14 185 -10 208
rect 10 186 14 208
rect 32 186 36 208
<< end >>
